// Code your design here
module ripple_carry_adder(input [07:0] a,input [07:0] b, input c_in, output [07:0] sum, output C_out);
  wire [06:0] c;
  fulladd a1(a[0],b[0],c_in,sum[0],c[0]);
  fulladd a2(a[1],b[1],c[0],sum[1],c[1]);
  fulladd a3(a[2],b[2],c[1],sum[2],c[2]);
  fulladd a4(a[3],b[3],c[2],sum[3],c[3]);
  fulladd a5(a[4],b[4],c[3],sum[4],c[4]);
  fulladd a6(a[5],b[5],c[4],sum[5],c[5]);
  fulladd a7(a[6],b[6],c[5],sum[6],c[6]);
  fulladd a8(a[7],b[7],c[6],sum[7],C_out);
endmodule
module fulladd(input a,input b,input c_in,output sum,output c_out);
  assign sum =(a^b^c_in);
  assign c_out=((a&b)|(b&c_in)|(a&c_in));
endmodule