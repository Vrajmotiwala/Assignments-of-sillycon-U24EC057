module ha(input A, input B, output C, output S);
  xor(S, A, B);
  and(C, A, B);
endmodule

module fa(input A, input B, input C_in, output C, output SUM);
  wire S1, C1, C2;

  ha h1(A, B, C1, S1);        
  ha h2(S1, C_in, C2, SUM);    
  or(C, C1, C2);               
endmodule
module multiplier(input [7:0] a, input [7:0] b, output [15:0] z);
  wire [7:0] p1,p2,p3,p4,p5,p6,p7,p8;
  wire [7:0] s1,s2,s3,s4,s5,s6,s7;
  wire [7:0] c1,c2,c3,c4,c5,c6,c7;
  and(p1[0],a[0],b[0]);
  and(p1[1],a[0],b[1]);
  and(p1[2],a[0],b[2]);
  and(p1[3],a[0],b[3]);
  and(p1[4],a[0],b[4]);
  and(p1[5],a[0],b[5]);
  and(p1[6],a[0],b[6]);
  and(p1[7],a[0],b[7]);
  
  and(p2[0],a[1],b[0]);
  and(p2[1],a[1],b[1]);
  and(p2[2],a[1],b[2]);
  and(p2[3],a[1],b[3]);
  and(p2[4],a[1],b[4]);
  and(p2[5],a[1],b[5]);
  and(p2[6],a[1],b[6]);
  and(p2[7],a[1],b[7]);
  
  and(p3[0],a[2],b[0]);
  and(p3[1],a[2],b[1]);
  and(p3[2],a[2],b[2]);
  and(p3[3],a[2],b[3]);
  and(p3[4],a[2],b[4]);
  and(p3[5],a[2],b[5]);
  and(p3[6],a[2],b[6]);
  and(p3[7],a[2],b[7]);
  
  and(p4[0],a[3],b[0]);
  and(p4[1],a[3],b[1]);
  and(p4[2],a[3],b[2]);
  and(p4[3],a[3],b[3]);
  and(p4[4],a[3],b[4]);
  and(p4[5],a[3],b[5]);
  and(p4[6],a[3],b[6]);
  and(p4[7],a[3],b[7]);
  
  and(p5[0],a[4],b[0]);
  and(p5[1],a[4],b[1]);
  and(p5[2],a[4],b[2]);
  and(p5[3],a[4],b[3]);
  and(p5[4],a[4],b[4]);
  and(p5[5],a[4],b[5]);
  and(p5[6],a[4],b[6]);
  and(p5[7],a[4],b[7]);
  
  and(p6[0],a[5],b[0]);
  and(p6[1],a[5],b[1]);
  and(p6[2],a[5],b[2]);
  and(p6[3],a[5],b[3]);
  and(p6[4],a[5],b[4]);
  and(p6[5],a[5],b[5]);
  and(p6[6],a[5],b[6]);
  and(p6[7],a[5],b[7]);
  
  and(p7[0],a[6],b[0]);
  and(p7[1],a[6],b[1]);
  and(p7[2],a[6],b[2]);
  and(p7[3],a[6],b[3]);
  and(p7[4],a[6],b[4]);
  and(p7[5],a[6],b[5]);
  and(p7[6],a[6],b[6]);
  and(p7[7],a[6],b[7]);
    
  and(p8[0],a[7],b[0]);
  and(p8[1],a[7],b[1]);
  and(p8[2],a[7],b[2]);
  and(p8[3],a[7],b[3]);
  and(p8[4],a[7],b[4]);
  and(p8[5],a[7],b[5]);
  and(p8[6],a[7],b[6]);
  and(p8[7],a[7],b[7]);
  
  assign z[0]=p1[0];
  ha h1(p1[1],p2[0],c1[0],s1[0]);
  fa f1(p1[2],p2[1],c1[0],c1[1],s1[1]);
  fa f2(p1[3],p2[2],c1[1],c1[2],s1[2]);
  fa f3(p1[4],p2[3],c1[2],c1[3],s1[3]);
  fa f4(p1[5],p2[4],c1[3],c1[4],s1[4]);
  fa f5(p1[6],p2[5],c1[4],c1[5],s1[5]);
  fa f6(p1[7],p2[6],c1[5],c1[6],s1[6]);
  ha h2(p2[7],c1[6],c1[7],s1[7]);
  
  assign z[1]=s1[0];
  
  ha h3(s1[1],p3[0],c2[0],s2[0]);
  fa f8(s1[2],p3[1],c2[0],c2[1],s2[1]);
  fa f9(s1[3],p3[2],c2[1],c2[2],s2[2]);
  fa f10(s1[4],p3[3],c2[2],c2[3],s2[3]);
  fa f11(s1[5],p3[4],c2[3],c2[4],s2[4]);
  fa f12(s1[6],p3[5],c2[4],c2[5],s2[5]);
  fa f13(s1[7],p3[6],c2[5],c2[6],s2[6]);
  fa f14(c1[7] ,p3[1] ,c2[6] ,c2[7] , s2[7]);
  
  assign z[2]=s2[0];
  
  // Stage 3
  ha h4(s2[1], p4[0], c3[0], s3[0]);
  fa f15(s2[2], p4[1], c3[0], c3[1], s3[1]);
  fa f16(s2[3], p4[2], c3[1], c3[2], s3[2]);
  fa f17(s2[4], p4[3], c3[2], c3[3], s3[3]);
  fa f18(s2[5], p4[4], c3[3], c3[4], s3[4]);
  fa f19(s2[6], p4[5], c3[4], c3[5], s3[5]);
  fa f20(s2[7], p4[6], c3[5], c3[6], s3[6]);
  fa f21(c2[7], p4[7], c3[6], c3[7], s3[7]);
  assign z[3] = s3[0];

  // Stage 4
  ha h5(s3[1], p5[0], c4[0], s4[0]);
  fa f22(s3[2], p5[1], c4[0], c4[1], s4[1]);
  fa f23(s3[3], p5[2], c4[1], c4[2], s4[2]);
  fa f24(s3[4], p5[3], c4[2], c4[3], s4[3]);
  fa f25(s3[5], p5[4], c4[3], c4[4], s4[4]);
  fa f26(s3[6], p5[5], c4[4], c4[5], s4[5]);
  fa f27(s3[7], p5[6], c4[5], c4[6], s4[6]);
  fa f28(c3[7], p5[7], c4[6], c4[7], s4[7]);
  assign z[4] = s4[0];

  // Stage 5
  ha h6(s4[1], p6[0], c5[0], s5[0]);
  fa f29(s4[2], p6[1], c5[0], c5[1], s5[1]);
  fa f30(s4[3], p6[2], c5[1], c5[2], s5[2]);
  fa f31(s4[4], p6[3], c5[2], c5[3], s5[3]);
  fa f32(s4[5], p6[4], c5[3], c5[4], s5[4]);
  fa f33(s4[6], p6[5], c5[4], c5[5], s5[5]);
  fa f34(s4[7], p6[6], c5[5], c5[6], s5[6]);
  fa f35(c4[7], p6[7], c5[6], c5[7], s5[7]);
  assign z[5] = s5[0];

  // Stage 6
  ha h7(s5[1], p7[0], c6[0], s6[0]);
  fa f36(s5[2], p7[1], c6[0], c6[1], s6[1]);
  fa f37(s5[3], p7[2], c6[1], c6[2], s6[2]);
  fa f38(s5[4], p7[3], c6[2], c6[3], s6[3]);
  fa f39(s5[5], p7[4], c6[3], c6[4], s6[4]);
  fa f40(s5[6], p7[5], c6[4], c6[5], s6[5]);
  fa f41(s5[7], p7[6], c6[5], c6[6], s6[6]);
  fa f42(c5[7], p7[7], c6[6], c6[7], s6[7]);
  assign z[6] = s6[0];

  // Stage 7
  ha h8(s6[1], p8[0], c7[0], s7[0]);
  fa f43(s6[2], p8[1], c7[0], c7[1], s7[1]);
  fa f44(s6[3], p8[2], c7[1], c7[2], s7[2]);
  fa f45(s6[4], p8[3], c7[2], c7[3], s7[3]);
  fa f46(s6[5], p8[4], c7[3], c7[4], s7[4]);
  fa f47(s6[6], p8[5], c7[4], c7[5], s7[5]);
  fa f48(s6[7], p8[6], c7[5], c7[6], s7[6]);
  fa f49(c6[7], p8[7], c7[6], c7[7], s7[7]);
  assign z[7] = s7[0];
  assign z[8] = s7[1];
  assign z[9] = s7[2];
  assign z[10] = s7[3];
  assign z[11] = s7[4];
  assign z[12] = s7[5];
  assign z[13] = s7[6];
  assign z[14] = s7[7];
  assign z[15] = c7[7];
endmodule

  
